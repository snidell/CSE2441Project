library verilog;
use verilog.vl_types.all;
entity Selector21 is
    port(
        Y               : out    vl_logic;
        B               : in     vl_logic;
        S               : in     vl_logic;
        A               : in     vl_logic
    );
end Selector21;
