library verilog;
use verilog.vl_types.all;
entity QuadSelector21_vlg_vec_tst is
end QuadSelector21_vlg_vec_tst;
