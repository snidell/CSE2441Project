library verilog;
use verilog.vl_types.all;
entity partA_vlg_vec_tst is
end partA_vlg_vec_tst;
