library verilog;
use verilog.vl_types.all;
entity Selector21_vlg_vec_tst is
end Selector21_vlg_vec_tst;
