library verilog;
use verilog.vl_types.all;
entity InstructionRegister_vlg_vec_tst is
end InstructionRegister_vlg_vec_tst;
