library verilog;
use verilog.vl_types.all;
entity accTest_vlg_vec_tst is
end accTest_vlg_vec_tst;
