library verilog;
use verilog.vl_types.all;
entity accControl_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        C7              : in     vl_logic;
        C8              : in     vl_logic;
        C9              : in     vl_logic;
        C42             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end accControl_vlg_check_tst;
