library verilog;
use verilog.vl_types.all;
entity overflowDetect_vlg_vec_tst is
end overflowDetect_vlg_vec_tst;
