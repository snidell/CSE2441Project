library verilog;
use verilog.vl_types.all;
entity accControl_vlg_vec_tst is
end accControl_vlg_vec_tst;
