library verilog;
use verilog.vl_types.all;
entity opCodeDecoder_vlg_vec_tst is
end opCodeDecoder_vlg_vec_tst;
