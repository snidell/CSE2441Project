library verilog;
use verilog.vl_types.all;
entity controllerTesting_vlg_vec_tst is
end controllerTesting_vlg_vec_tst;
