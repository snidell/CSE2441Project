library verilog;
use verilog.vl_types.all;
entity FlagRegister_vlg_vec_tst is
end FlagRegister_vlg_vec_tst;
