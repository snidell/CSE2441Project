library verilog;
use verilog.vl_types.all;
entity addersubovr_vlg_vec_tst is
end addersubovr_vlg_vec_tst;
