library verilog;
use verilog.vl_types.all;
entity controllerTesting_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        C1              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        C5              : in     vl_logic;
        C6              : in     vl_logic;
        C7              : in     vl_logic;
        C8              : in     vl_logic;
        C9              : in     vl_logic;
        C10             : in     vl_logic;
        C11             : in     vl_logic;
        C42             : in     vl_logic;
        Jump            : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end controllerTesting_vlg_check_tst;
