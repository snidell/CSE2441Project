library verilog;
use verilog.vl_types.all;
entity partA_vlg_check_tst is
    port(
        C0              : in     vl_logic;
        C2              : in     vl_logic;
        C3              : in     vl_logic;
        C4              : in     vl_logic;
        C7              : in     vl_logic;
        C8              : in     vl_logic;
        C9              : in     vl_logic;
        C42             : in     vl_logic;
        IR0             : in     vl_logic;
        IR1             : in     vl_logic;
        IR2             : in     vl_logic;
        IR3             : in     vl_logic;
        MAR0            : in     vl_logic;
        MAR1            : in     vl_logic;
        MAR2            : in     vl_logic;
        MAR3            : in     vl_logic;
        MARHex0         : in     vl_logic;
        MARHex1         : in     vl_logic;
        MARHex2         : in     vl_logic;
        MARHex3         : in     vl_logic;
        MARHex4         : in     vl_logic;
        MARHex5         : in     vl_logic;
        MARHex6         : in     vl_logic;
        MDIn0           : in     vl_logic;
        MDIn1           : in     vl_logic;
        MDIn2           : in     vl_logic;
        MDIn3           : in     vl_logic;
        MDinHex0        : in     vl_logic;
        MDinHex1        : in     vl_logic;
        MDinHex2        : in     vl_logic;
        MDinHex3        : in     vl_logic;
        MDinHex4        : in     vl_logic;
        MDinHex5        : in     vl_logic;
        MDinHex6        : in     vl_logic;
        MDoutHex0       : in     vl_logic;
        MDoutHex1       : in     vl_logic;
        MDoutHex2       : in     vl_logic;
        MDoutHex3       : in     vl_logic;
        MDoutHex4       : in     vl_logic;
        MDoutHex5       : in     vl_logic;
        MDoutHex6       : in     vl_logic;
        Mout0           : in     vl_logic;
        Mout1           : in     vl_logic;
        Mout2           : in     vl_logic;
        Mout3           : in     vl_logic;
        PC0             : in     vl_logic;
        PC1             : in     vl_logic;
        PC2             : in     vl_logic;
        PC3             : in     vl_logic;
        sampler_rx      : in     vl_logic
    );
end partA_vlg_check_tst;
